
module tb_FactorialCoreTop;

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "ModelSim" , encrypt_agent_info = "10.5b"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ETwxordrQKZMKw0YESTsUO7lNkO9QCQpizmHjqyFOwI0hSAkjgUePxf69AUv44bq
avZX4G/YMDObClQt5GsNcKraUZ2A77MphDfAi4RKzZCh7TXlQ2O7H+hq9Nzjar3T
p+2sxZKydw/80/ZIZiXaFU3b6hcFtIpZ/H0VqN9eFhUdKgJH8bpXKnKmXf/dEqtQ
I/Wa+OgcH8yhVpCs5T/5bs2n/ocJ9wJPwu1eJXKN0p/OhRiHPevPklM3JclFKKUH
cV2OtDqC6utaSMDpiXpb2wuSjGbB/yxMqDSZUMweSQCBme8MXaF6iWNRZ/jzdDj3
5skdQuv5DbM3HDzGG7CHvQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9920 )
`pragma protect data_block
WiQfTt+fW+LrCuLFxI5+1K6XZUtTp+GA9RwMts6qy2i3XCEVYZjvQ6Ff0WaxkfEy
ztSIQ0diMn7SC+N49GZJZarsOl5+/iqj9HbEQQfSfSVZ6JkszKbkQ1FLOSpT0KtQ
jbY5NHexHYs2Pgvd6qE9bf5uTEtdzCpAud9vYBqR+e5eWjpLHfiFFtfSxEBKBWiC
R06HCrYoNljjrczj9AK8hAISQ2iz1uOP2WzSU7mNcAw9pmQXzllYTU1Rw06SsUk+
oJMpPpg1bDxtOp3AhLP+34c2ZDbzc4j4KpXCINyP9OSVxx0a1TdxjJHsWtk8SvSY
C6WNbGgLvoH/otSFJ7OZgzCkqO16nb5iCoDIk1wfKdK328y47Q4vFClE0Ar8r/0m
i/LF10khECb0byHdK6x1zvmaGWt7zJd+NvpWl6kT5ZcA3f/TZyVB8UeZ0MSJmbhR
RE5gm1nlgQKRZImEkuk76D9w3geRISVwfHzGDIUMJI/iDSDTxQZQ2lhDgwC6kKDx
rAu7hTTBWGNYI/sR8/lai2J/P71dhtwSMJkzOV1GS0wBCSPHT12QvxmqmmKFZEKg
vcb70AC6i+j1pNyhvepDrJ/C39Qq6TyHGuBah1Wxlt82Oj633LYsycpvcHBJMCfj
F1S1pwfjVohrkH9TGvGHn7oOJSHLSNEHfRY/SI9CNtz/Jj9e7rvzOuruebRE6nry
xQ1em38xc98TZPEdDNg6HwOvzyIQJvQw5qfkJCNFcq2W0aeylwCu51pn97JjKUGD
qlGi2lQmK9qpPG2ifQQ7gDdbH19oFmPREnTpqFYyKshvBnoV6qh7peRjZvvyP6Lp
S8k2d3WjL2ZmFdg4dfk8/NQlCZQ47iYAvOzl/20ihARNOoLZBaP8r3P5ypk0xg2P
4RmhECBBRm1nQCxrJ1Y2P94q7FmfgxeJbc7bCkBxaSC3StlpBEz9EOaNVA8QT9Ve
LGD9qYUnRCpyFLxc3UKU6AsLm4bmgJPCPZmRx3wUEtwgne7hNLPC+TTQ1xn7UKyj
Wzyp+iLQXOa/vO0ptoO0+6Teud7VqP1Vt+cuEAzInkWccSZay0RbwL8KU98w0KIE
WzDY3LKuxQs+Kc4xnHVizz52iwtA+0s5DlOUSzvI52dJhNkRQPgeSmY7/ROGBfEZ
rnmbKh10QL2aXvPK0ViwWFAv0qmVUR5HY/S7pmXr1PtdQo++eWArKIPj25g1EbMo
G2sQXuq79IkfGFIbWkPQYABDk0GmmNm+4JgcvfWdJyHgIlOoMuw1JPYaTpGBFzRN
6ULnT7bAVLj3VguvVERgRjXku4pqD4PEUsVeqFm5PukXeWS6mxEeMDSAA0lRcIC2
dfrsEr6zssZnjZIcbJIE261WXrKt5mBxY35gRQAa52hwwp6I/nPzDyEjCJym79D8
p7pjdqRDMhJOIzTvyE3yAFnZf++y734DqXtKvVfM76UizxOQy7pZ2B09+zd5dezt
Htj1HlJCgYbkd7C2V/jRtY3MY0QBXMg5MZA9nXLQ2f+5aVdzz2ZOPFBy1lNF/pr+
zDBRYSqzhXX3IISvVNNF/3zOclzKc5G668NTrgONMGhFgcQjZYq31boaMJYSIq38
a5p8Af9oquS0Danc8U6TBw18Jat/za5XVUCiCsmI7FDxIVn7rwEhvlDdgj+6eRrM
S1aBkQDUm0SQCvwHsxOJh9s0OLehdisPec3YCW7OnAbUZgj1fYzeYLV3FDirLk3c
cMfCz6aRjZlP95k4gSJPD6jBjUfSiQlFMMSRFHy93YvaT1vzEFQZUOlocsAXkRbU
2lodVZ2BU1FIz8BolzdFXHxzwmZ13novMd9yykaEhJJ3oiGCtUadPCZrQlenJ9Wd
48ZFkogMS/MJqUMvvtg2p58UGP8DBAyo3bGsb/4YQ20zfbTtOp6pZXt8GCUcmBdF
Jf1i6oBlN+XsWGLfpu7ViBvRBsH2PSAttnEWlwI9qz5WqfCxsycdu0MJpRxDSuBg
fruwDPc8qOLaQZI/UMDBWrZakgPiXgQf5nf3G3OZZ/NcYWcpRSxezdr5Vj4px8i8
s0idCx2qdGBNNtrgevh/wsqnw2Os9Zwlr3F6weKNCTZiqMCWa8tr6IWNl6LF0JRx
+Wpqc2+oOUsnFLPwGjqCO4as57HumdxN5B30NizJDZYypT+sqN+RmsW8ORbi3+oF
qCnwvizbm+cFZ8ArPzdkI2c3VBnP6MKnsN2eG4tzeQA+O0c+hM8MbyDRUM5RYuE/
CaB+T2VF9mKioDdUjZKXm9EgXUWMydAE8GdOniS1YE28/ZaFWdXQT1yr1QF14UZT
3LuBt7hLTNewwTKzqexi9a8cHkS/BU91ZJ3g3zKDt94qWM+wNi9hCBkYWDlrVxMa
rkdDbuEd/W5MCOKiUIuM61SFDENX6y5CskEppjlLhzHxZxAx/3dvA3C8pXQNxeBZ
sxVbv75sEYWaGhEakSlEmSXAK8CAAOWj0WrqhQ4aFQCte2GxjiecfxdcFyfglczY
ZtBCc+YWO7sEDMxRctTGE24zKb6ajW8xycnSfXS+rUQ927Cm+aWHxobrRidH21f7
VGcwLm/HTAZ96EF80zMWNWDt9KQcJsyAIh4hjtUiiI86a79jpK5+/6zXFW91bSny
rXSViHuPn8xnrLxOpAQy28hDn/ID4ZhIYhjydtkFwraPDRAANKbFzRAc13S22pvF
I8y1wornL5TLekTXGbHOj/xOVdElrObIIR3gRdMk2vcQMAsKpCKxRJPtM8PWzHGr
5vCj0DHfyCe8Cn7qwx5Mzi9ev83d3mO9BUaz1LbDlr6kFueX8Uv6ZpFc5hGAa8eA
CLvYLcQy2EiU4WOjb2ayFPqtuIhSMsq+kO4AliX+AWcK7BsyNb0j7k6K4WV/LdoY
NaJlipNhQ3cRtsEUe4bFpbjZ4/8plzRcamud4Q3vcqia8IC3oIxWpjQvOLhmOLgb
29VIm1lUHJQAH20gHeKOfx10sVOIEgvPZwTuOZaf0zvAKLgCqAqkzMdEuwqozh7Y
eYC1zYVZ0k9kb6k5HQe2ZUc2F/xnKg8SCFayoK3WyIn8rQ57gI54hrwNO5dBXmQd
amJNCcCjzUZ62LvOJiz0mxcH9/nLXcSKcRqM2IG93pp38sTnuSOv+ei8mQJCZ1LC
YIyCmtO0J7zu2QkZlgbOvMcEYbcAal1XBOz+uAHQu/z/skhK7uxTwNXVGAZ7VbaR
7gECOvTkU3cyTWPg0eoClpwnyGgRytQIU7QY/qyLu8+U+mwOCSii5pFu5YeU92bJ
dLsaFIGMFvD1j7hLLSvKAP4sAL1UdJKvqa6vViF7M2AfvC/M9Ks84V+xdHGzxpqm
bITdKCU6txQzWs5ud7ukivwS9w9A9LOOpD9G7d3tI3ylPYwq8cb/NAApAgDQgxpz
/Ex53rYXFYPbgEwVZPvFlesk+5MvT/EByJ8POAWyjLzq1cn/KkKO9RZ+acnJsRec
b5Sgka3Pa8Ncq+RgZSkqwpgaVURIESnZzoSyo8gzIjE1Nlh71OobOGZo809yF+cY
oDffNUAKDywuBiMjXk8Pbyz1v8ZKF3Mehnov0ZEUzLG2J903Ez7eQ1SV8f8ttsj0
+V1zhky+L6jnVgoZMussbyf93z0VsxR1qLbkoxW/klmnhpkJDw4Fl15XAeCb4uNl
1Nq2CJoRq6V3EHCkJFWuRWGidud+JlmshqLGYjhtHFsysJlBRK4IcwAOhD5jr2Km
KcJj4NjBGtHUe7m3icrgTEF9tR6DadB9ccPOIdF1mf+WHi/DqbsW2LS+1CRGuKTK
VEU7AsyUX9jDqOOsSCBqRD9U7THaGk0gYHe0yJLuhOCRPoW11HpunhXYVYR/Q5N6
10K2FH+gkb1tH+lO3Ho2Ns9JA0InoETM0dV2e+k6dBljVIipK2ty+b41FhdLWjPl
JaMk+VAPfTTSH+MCftY4X1rRAdqEP1iIuGL22NKgnvKmYn5JJucb7SdvZ5cqu+yc
NOAhSEU/eohDb9ye/t1Poa9LOQLlmnPiYnXMu5EY3qLsHAa1P5Nxweb7c7kSgdfq
wfPHrxUkQfbN2wHDs6pQJObBTHm5U27FDM3ZhiSxkL6quOjr2oPHSSeBl2nFwb1R
cDSPHc2X4uDEDppqkUb2HxnVXkwE0O7e4xqWs8yv6WVFRAuoJAOEpfJrGnjbzAqs
Rwg7ao7/xyXmuQxQ73BPhntaxpg59/jeqBXvDz2cXcDIzvaaXP3PpLTDaJCdta4y
ddUziCreHynfLTO7zwHYDPg+j6K9eGJrwlILT0galw/ie741raaCKpCSGIjIBQFS
wu5IYCXq/q4e4rmeylsTtdRwkBXjN90jDR4Yye87vpIGbwSfylebMZLH3+GPyQi3
6fiDSv00np5ERLXVDZLWPRQXRIb+6k2wjcHHA+lpeskPscsGYFJ1b7n7WULUIzCy
FZsG4LCK7q2PYDE8F1G0YyW2mdiTVQn4Q5j8BCbXVxCBcqa1kg9KrEl+QNR03YJ5
+lqcPLcZ+U2H4gFBlqVSX0ynDbtV8xGMox91WDMfwvEq0AUZlwvyTWAbpl+sciRq
6lLQkyzK9XWmJekFT8a7xWyBxQ2PkKwjehiZ2R/9G6kIe1EavOMaXIDecxE2VRl0
/rVt2o4BR97ADA1Qc7OlOlwDdTquoGHS4avkKIt+Nsrr29CIwYD/uFM0OdzR9+vd
/kz5QXmlOVWkBmYoIcdCt8VRAiZQlXGJHxGRM3GINHZivaZXTsXOgC0NggxYgM00
Bwgst+GMQ3iQ0fgjDRzcBr+KihFSHj0MUd2fFd9/yaky06lviIsEw/IeXYqOfLCQ
eTXcPOjB+ybC8skS33E2Eji4Rk94220YbG8NF/0c23kRyDReXBM4eMAY5c3rfy66
2RBTRyaBkHDLBDS4l+TkBb0K/b5C0947hABD875v6s78Sk/p0FCv1WCbYJo+ox/e
d0hKqggZczTs6E054viw+3gsXzagPKNB3fxZuxmEW3FG2yrzR4Jl/vwJP00zPhKJ
Wco/iKVEQjEq1jvSmM7ODsBeHASc4o288fDtfPYnpCHqf6nNIJtsEQzenTfBhTuS
rmzv8woM0hP1frMCojRUAesioYKXU2hRaw9+Gx9dI6b5WUrnEgWZJJoopPaHW3mx
wdw4r6a0PC2kDYrUqcS8GqkPsR00fYmLrNDUcodrfCTkRk4Q16FuFTtY54OrArsc
rdGjdN1me4U7gSfcYYWWd1crA7yq85lnn3NsL2UMzl5prhz3amfhpArjnqxCpf5m
m/D18wP17os0oTJ4dd5w6/5IHjmzobQQnM2F/mSAxOCiIEGlq497xIdnJlLVzSAb
ka4QjPOCEqfRj1PiWgxyQvKrAVLet/yLwxHbvNCtDu4Q0I0xfDfyOcQqDCjaUFw9
GThlQY1pJNKZ/PLjyR1tIhvdeqnyZcqG76BhRBGLmy4vqDCv3vKC2pRNTIZi+nIX
Vdvi6gTDqbudftRig3BbFXqSfpWOHoE8c4kIqBVSuuAh1ySPGwqP6Z54ZshdLo8h
EPI74rYME0pyTWXwbxf/C8ZDtlrefRl6gCr9Gk4vgTEXbK2gLIFqKgQcO4ziJjEA
Tk2busqBFLs+7A+QzDAMuy8Qer6OwKemoXICzCzqzT2F5gT9re4SahgvWRkUg+Ai
Xt8n9qsHKdMKGWoTLimRhQ3pfJz0bo8vloTFuGktfW2uFwPJDUqLGZLT3SmyCpxJ
q1URV59BDjwHZpVgxLC2gTRlat7UHXcB+v71/9Yg/rbTaVfEAKVmgeKcKwDYJhLl
mHf0E0wP87fIiwGWrytCkI5Zswqe/EAn4HjoFd8+SxjkuVAOdIoCSqOcmSjd5WDa
eqsZ0Da/x0Dq2lfrgoD3n0a/17lnmu0saWyaLUs38jCL9OM1oPND3o2/q8jDqe+F
rUEOC2y5H8IoYSkfPldPYfeF9EhMYrW+VBNTnf93dyiXcXjdyxnYC/1XEnZMU3Mu
iXSgh+GHd6G1nju+y/CXfehPzLeKJYD16CDLtx6fGUNxJC6b79PaU4QgLHwzPNP3
iEVv3a/on2PnUVyXVxxNmO5qrrlIt1i4/bbLBBX6wwkQ6wkercApzokK2qSJitnz
sTPxxG0++5rIcNIswRsaGoq/tUKifU0vC6jGCPKVuwZSlA6B5DqccfDQ0hZ9CFMJ
27upwnfdw3dNE/it28h6/k1HYBdAS9RKQj31UM3H3UnpTBKb8U3TB0wu0tnWbYkc
0aJwOGGor1xJ4jM6QPW5RPe8593Rt1Ob/U3nJ0B+GUYsdeq2Fwzi+udpcQtBPclZ
aV1A57Z5sH3WT80BnGYTtgNCbXc0EJpQD0e/0omce3f0nrLySUL44QHdLKhaIIe7
HZmx2COXMoj04Y5q06glqbn4wmbZAiXy8a59Cf2wA+9iG8X1lNjFu1//xLX8k1X5
NGXnLtq0uTiDyG1pxCpA8AnGTKD3JGAkE9+3FdYMPScPtaa7tdo3vM8tNziDOG3y
Mb/NS1+E1jG98xH03m8XRkvpyMBJizT0XMsqWbBan2V6fVzwsoOkdtrQWX9ZmN0I
nzxAZmFb5DCtjlWeWE0fZetGbk+W264ywjhn+81fLOELeV2QNyApwHPkLRHYDVd2
XXvbPwwtCjCrGYf+HyF2A62O08y7UWFoI4kfjkihdtKjfudvXiF0lfNAWnSLcVyW
ZzYl0u904Kgf/qebQzjkO47TWUN/YGYlTzWJwoBpJe1YsaCrqW4nY3rMRo9riln9
eld4q6DQa8WC/AQ7bjRRcNCaOSm/EZPJ0N8THFLFhA57z7pErpiFGE2UXnnXuozc
dU8Zl1oAc9qT7lQvifV7L2FcaW0h1CQMVJC1hY0Urxu2DBE0MmXcvMgL9xzBe59b
hPun+3NUYZoWsfYl4A/iEQxnsd83KSV1fX+yxQZ7VixD50+pKffV5xIg6oUnPAkW
h1N5/QH1aH6HcBRjqGQTvyIBLBaSUQYFCxy2nH5/sjcFJhgs4oFEw1hCJSQaxj7y
SNw5gBcdmJfcabX8whlvxHSuc3Sn+jllAZMUSg3MvhDx2kEpL7kYuJE/6mcEl48e
6JZtgOeNBs3dB45al7RcoUVzoUuDhRy4lwE/xX6F4avlNMjrVcvv2INXcjAPvB/s
zlSAWrWADDlrP7stCccfxf0A+xaBys2Bmpa8qSfrIWcOFhI+q+BdQuy+R7SWyq2V
SUv60wofbbqbKJV0WR4DNcrkrZZULB0EyKFBJBrct48C99rDX9sMmuG+8rL1iY4B
dHjG98kY2geJs2C3CxfbwzwKUr+8hD8j3YsR+YMPjPJRiXG0PGKDJCjuEld0Q9+v
IXKtB1KCQ8GuhCwaXZOD0nzGZMnVCyy6CJl2iERsLfloY2CADlEVK8+N5f2xYpnQ
22ueTb7Zum5nlTSoWu31z6O7FebDuIa0k/FbLRQfntYkwj7jHHmxOMKicVDj6G0E
+v2RgqPOkqqZvoLIvjyTb6MGhc6x2ecHFopi7ns8wefUTtHjZWEDAhJp2hK4FldR
f7Dm1koJxDMxCxzNuyckCLn9Wyeizn3U9Bdx4sPzovoCS/iGg6HA++2UIk9knJu6
Z/osrizBAkI7WyaLFctgtX2DAfNVCEpYYymFiIepZB3QSuvxFIcdHPOMN4so0vl2
9ste52tvcFGXs7OvAAO2uUwG1faBubiVmIIVI7+wd6ha0Zfn3QIB5+eqWci68kPX
xYMb7bVFmuOQB6YD2A2F8kbbeKUep70nIbKeUfJp2s+6Q++EOw6XRp0Lj9PzwDqA
Ql8LFXlyvxMWBeU0nrMt5gXgScL1FBu2qDCTQPXUIvVnXCZq8XY/DPSvkQOyCXjy
MmvFihKlsj+uxnF+gUZAYTXGiunCQT/O+NzffuooNmKjBBK0gxdCKseul2hXhr4i
6OZZ5K9gVu7j+Fz5V7SWih3crjkOJABNKhHmizV8rAqgkDbLIsadRQ/yspDTWZ7W
JO0Klx3k0jRlZfYV5/G5xQunOviCf2Rktl6Ta+xzlExXNM0rSL3UgijvDB4JLz2p
svIxJ7u3FZiglJJCyqQvquua1PpbxSeJ7M76Pu5w/twOuw39dAcUWF+dEslWxCZc
HwORyW+orVkp7JOL/M2zo9wkfaVEHXHYqiu5bs2iFupJyXrp/hGanspY7pHySoiG
+TtdSG5Z0mCwLI2tcJHX0fzaHpD7A7GYRYdtHLiMsWfnG+WNiVbTBexHn6RnQNuS
BYiKVljO8ZGmg9AXMQz7myZJAwLYQBcoAgDKGo2wyslEK3bGg3K+whDxRAC1wmV4
AUptwAfPafgTlmOfneRQupcNlDH1UpEHBgIDcg+myJYvUgnMRXtgSzA4p8OgW+pg
/gK/A2bzBIUP1WquOTk1CFAUkLt9hJ56wnyeYjMiUWkABHinIMX4asj10MW7+/S9
21gBYBBMwWA+EFslQSh0pNKhGqMRUM4mHB+uqyC8jdL8tluBbMIuk6ob3C9er45V
UCpkKCrm6KyIv+xRiULPYR6K+pfzmiY5KXzMdrpou+Q8SeTcFxtBMMwhD7rq1Of0
WPzKmHnEyVYyvmdDSotCG7lWpckn2aeuJO0Pffcumyg9P7P8GRDrvhiV5xYCllgz
aA1kZDcaOEMX0AYIIKgQ+xZdXHiQ3WrHiBugIA40uyi1ZC4l1xnX+LFHnNr9FBT3
vJV3J1V7yN15en1l48a3ueRJ5JQkPPXc3RTXCaKNr+AjxVKlXRXOq3TM/cpkuFuz
aidXmPwfRWqFekmkpHPnJDcMJ3PMM03fAj6PF/JZ8nShhRpyccRTlzvKLdyfw5sr
yGWPzVTq5lsl2pl2iVfeil3qLNBUHXyN53y7mR+Qm9TxN6nNSQtR2Lgg0pklWNvS
27TMvSjAZpR90cjDbEX0iE1DvUkLjc/5Bg1BWEvHAe8oaPosgop7ANtRJ2vQeisj
0G56idPYXI9lQcFbdF/eG/7HEcrY0Z3ViTYiHqZZP9rW3bdAbzlvuBMsmRVYWFKI
XPWM+SrSEqj5+JOcLQGOXV3XSfbOrvlwP3XJ0aA10ttaj032awYv0TmZnOlbU1+9
GFoFt2XTyRSFLnCUr49jd0CbM7Acv4vYKDRFDkxqQZ3H+/hHILKm0sRbvtp/abf9
pz2S9kUU4QiGNdwheLwYoTf602gzgQXw4ZKsBOowwtiN+hOLUa11xeFldYgfYJRV
CheBU8RQ1SOhp+Cpho16IJybs6jQM6p7lC4vTuU7LyCbjihmzpEcTr/VGMkwQdT3
XYUzE0tN3e6vBeuZjTN6fVv1u4GcvXdljipTKkO6aG+OjHJN4l8uIao6NQb/U1Iq
6PBl4PVIlWu43KmyN01YFkP5j9vpmfXSsqUmhtqmlMTxfJmJm60qFTBSf8r6LyKY
nbN2TYl3TmxWi2hMOnlG//yZt10VE7y28eEHheBayujhtpilSOTjUPuGFGm9SYhs
ez3Vg3LScYRI7o9ag8pSF3FpSLJaxWlNNHbAhqmnhh7M6nBHHl7L5B5BVSlLQlBr
GLJsx1OsiHTZ9ONYxEZ8ssaEAoxs8Bb9DlR0V8Y4lC6DIgVnhIrqyhwOFuKETDQ5
SLyrC7RliuJMKUJMY7whYLkc5g9uBZ4MEvh1lBBeaQJ2Vkg/npAuWcUoj58DVB1f
Ugvl0tlXP9l2SOuOOc2prPP/Cy/JXqICUior8HYWiZFBiWbBRdhLdfOI56E4TBNd
13XEVBe3bgxPf7Vu8SAoVuIKR5/5N51gR0JIA32dmqKNIZPGoZHR9jmm/O0e/7hV
UK8Qd+wLeDaRhr9lZycdB2yacr6mNphkM7WhBvjAA8k+Zk9Z0zDn6r5/k9KOt/xt
FEwfm4wlQvwfYTEPXmeGHkWTnnmNPGp6vgPZXDxjSiQ0WP+L7DFk2gMhG8QknuwR
NIPyMi7aR+92jwAm6DIADPRsF7YPhwyaIfFwHg62feVxeUN1MhW0Lz6NU93ABC8b
+wRdckFv70VjxbLQDfCP1QmjpjxAe4jiXBtmNOJRjd630N5YrTbCqgqS793tRmdR
WxjrSNhjp1Tk8tLth+IMR3q6ToTVmsMkQISInFo49SQDCO9xooXwH4w3iwGQ7jiB
man38ixsKB0v73sIjWVBKrhp28mI5ZuUZ9JC9SJitfDL/7j5uAzLYu9zY40w1141
eferAoOodbA/Txri4EweWS1g5kugOUU2rOT0a7xuZSeo3t5t2xRl9z6PnI1GcOlI
5uILVZh7/Q95G5/jOhoyjkapJ9TXKJIZ6g1AVd5uXLb7W9qCW+loSfxgBHR/UV3b
K+y4Bgo97uVps0c2DtDYBfRQjbBJEF8cS45VBT1lXVN1bQJWOFCGW4Pl6DcLoK5Z
S71I+oBntpTAkyiIRUGpPS+twfpEG5uZ3D1Y3uIWw0mkKKkokq06VkrpY2dIYi+m
x27icFPkcjLX4dEHjmFf23m/uFhRD/3E0PEnYpLWEBPuE4ZVp44Ctejf19GIQX3L
jfvhtLzCwwHRwkdufmkWWN/11lT2oClD+HCIltCFUwJCTy4bKv099aYXc7pzXNl7
hgQj0a4xgq7pzK8uybCU/LvZYpqIcJkWmsP+etXtYEweVJkFBkQLkhhNXISLcUNp
XpCs3mY9uCdeWHu17NT765JrCMUueGUJjk/Url/X9gRDkjGPgG3b2+sUCMfM0ZoG
+37+prVYvY3bktiZnsyjKR8A5zyQ5NDp+cXLIIiONl0XeZKznXzCUlZ/u4tGnG28
Eg+NHb7PIr+r+JoZcL/l0gzAcOORJN/h/yDvnzspqqidO+3hflCKzbdkn57tSQaX
J/49n0nC4KfGdp0i+Z3fNbJH2jWzJXMKo0Yiz5Xupreoe5AkbXLS6O2iTK+dlTZ9
0njELxaJul+y5yY5EJwIPAuc6KZk1DRIMPtgXgc6OdEHWD+QoZeiHN7RfI3HQPfq
fXh3pWA30bCdKUqJQFNSiM56AHAF51W6zsdxoeMing9xERd9MpQG58AAAbbc5Qb2
wGwT1P59t54214YBVag4ms3ZosW3hqX0EDYYyeS9btlpoQYtskxguluca6NeIWlg
LSWe7kgKQ4LlsrBU9YXLaowzEP0UcVYyJWUaqQ9J8q0yu5oVLL+9PRtwRrt8AbW/
o0jrgN62BB3weaYlnK/S7PZ08noI2Zbb4MqQBuP2J/WduyttfJ1qi+DwsexyHwJq
a3bWP/jEd/rr8KVYkaNMz++MWD5m5BQQI4cAPxoCL/LNmKTMt5iDlQXFFw7sFNbM
r4mESlvnTNmW11YwBoGNfCDX067rZMKTXOtl2UYrk7zcako9rBsP6t28suKOU+SL
V8re8fWccArI7ojJIfL2k10es+kSDs8iYyaMTpzAlKWnFkowgDVjlbCH9hLgWLHy
lnOGu3nIOc8OJvU/InsjC8765ePsuxonrdj4a3rjHQuUkdpP7tyg4KaVNYmfwsKJ
4whTOjVDwGagX0Lru0eSjYSxLR2+AFiE9edMBdz/E1FCdfm3itVGoZNtXwzvwMqa
AEQhS7hzWu/jq7YKCJcHE2XZV9K15OiQ9WgG/tyzZEicBNUcA7/VuynpDEVa6ke0
fPRmfDqJox781xyWMJb2twwv39tyAEOkvkq8rMeV0E+dqCipJD5vhi7i+Ysk5svw
xeae3BAz2d2Ps2VYQQu4ERoManfR45IcsEebojHAPDISHq4fJhAwawaGHehRTaZ5
8XYKFR9K1EL3e+n1d05BGE+GGBwnSOAZFEstC8iUV+f2QheghDxyxaIemUeuXD8G
KdKts98dRnc235m0/YFJvf2h2M+vxTpQpvZIPV2rHGNXYA97iW0Ry0AvYC7FU/dm
Ffx+8U1OjCfGK39I2zRqYLSqUdifC8wTt1lA9YPegx90oFY0HfvBzOPmlQscjfs0
GFWRkHxsoVnFNv1R/tUCEkrwvMUiX4+ZysUOgxKSEC1PKz8cu4AsQLa0AdRLmuqp
o0QfxbVit1h+Z8YngRhCFSOxqwSj+fU0k3DmzYzExSA26Icra5uO+cVVB/Jk6e95
bo3g7ygjFxgwp0rST0F5jlpxlCzAJgjSgda6ZPXRvndbGxDYYJipQxJDqj/+6yr/
4IOexUnWjtvAuNt7ka6FvPUGgC9gB+WAes8Z4NzMEG1SWGwIeLQCBqNNI5X/sjjW
Qn18Ro7IhLI7vKrHo2oVRPcXkvK2V7W+5cqFN/pwiEBPNzi7xmaT2Z7iFBJiLkmv
cCqj1ICIrB5G5wnNMsNlk+ocrlRVISBVjEmH6EIDInxbhwgeAQCq8zfiTpTON8Ym
PqeHbjQQIxFk5POmqWy63zS3cUen5RZDrwe6EFOAVkUFR5FzL1EOsKOPMCRrjzkC
WIhjQ62tNFb6s9wypuVploSct8cEK/Ufpay5TmmElZIMTpALDtWPOp+WSO/fvXDB
4cF84BT+FV0fjBxnVidkwj8cXpb7fPlsgwmcv7qdPCwaH5cYd0IoKtpsLjMskYER
c53Ng1DxM3DrkVLOQLhzc25fR0VjK3DsbDLqtYhAnGhKOadnf2THM8W2AZu4kBCG
zLp1YtUukZ/Y2H/D1wNSdEewQKpu9HTc4k0LKgDnHhy9d0pRwi7A2fa3NK2gLH0+
CICgbPInALJGb4lpDO4h9dfaL4znF5LbAcnInFzjVSh6SI2riQwVpEZWFMtSQyel
sBbk94XzMutrc/DYzCkI/9PlkIY1H80HkOqR3Spun9Eq8I9crn1G54JHJSElBNMg
1RSMWCaxG0JZskCf0YtnNXWMFKUGwOzsnApSQJePM0jR3pcQV9bjWC/Ra+wD2uWm
VEBe4G4nEQaWo9fUkplhIbHUZ12b/N5UVx3PKNBiBJnSq5SEduUK4TT83gK2lz1w
oqnObJRenysYQCivmVXV1NWtnZiTOLSAwl1uqIthqo1Qy+Tm9Nyq8vbyv4n7URZG
tUBz2M90B2Upymkzt6jGQ6gJ1xtCaiGNAE93cszpjVrITsJkmFIGG77hpHlQHven
zKHg8Evow4YmqxnHtynYASup7/ovLULLv37ab3ah+CUazttJ80Q4cQgy03+l26sJ
FVTJPwbG0H33YcaJzvC5c1FajERgKDF92D7btaQF2mQjHo3sBCMuoikQOywDMjB/
NNuozEwwog+Vwf2k14cuohDe4bpugzIoNZd9wnmWOBOZD523qx3TaM0oAC11yz9J
J+vlImO4wadakWu/xD+LqSluXsrYX9yHikG909ujplmA3pdulB5ZBs8qHdb/mm03
aoNvAf2WovHPmgm/1kREWo46Pp359Z7ne6Fi2teGqqw=
`pragma protect end_protected

endmodule